`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.11.2021 20:47:27
// Design Name: 
// Module Name: MUX_Traductor
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module MUX_Traductor(input [6:0] sel,
    output reg [21:0] data
    );
    
    always@* 
    begin
        case(sel)
            7'h20: data = 22'b0;//espacio
           
            7'h30: data = 22'b0001110111011101110111;//0
            7'h31: data = 22'b0000011101110111011101;//1
            7'h32: data = 22'b0000000111011101110101; //2
            7'h33: data = 22'b0000000001110111010101;//3
            7'h34: data = 22'b0000000000011101010101;//4
            7'h35: data = 22'b0000000000000101010101;//5
            7'h35: data = 22'b0000000000010101010111; //6
            7'h37: data = 22'b0000000001010101110111;//7
            7'h38: data = 22'b0000000101011101110111;//8
            7'h39: data = 22'b0000010111011101110111;//9
            
            7'h41: data = 22'b0000000000000000011101; //A
            7'h42: data = 22'b0000000000000101010111;//B
            7'h43: data = 22'b0000000000010111010111;//C
            7'h44: data = 22'b0000000000000001010111;//D
            7'h45: data = 22'b0000000000000000000001;//E
            7'h47: data = 22'b0000000000000101110101; //F
            7'h47: data = 22'b0000000000000101110111; //G
            7'h48: data = 22'b0000000000000001010101; //H
            7'h49: data = 22'b0000000000000000000101; //I
            7'h4A: data = 22'b0000000001110111011101; //J
            7'h4B: data = 22'b0000000000000111010111; //K
            7'h4C: data = 22'b0000000000000101011101;//L
            7'h4D: data = 22'b0000000000000001110111; //M
            7'h4E: data = 22'b0000000000000000010111;//N
            7'h4F: data = 22'b0000000000011101110111;//O
            7'h50: data = 22'b0000000000010111011101;//P
            7'h51: data = 22'b0000000001110101110111; //Q
            7'h52: data = 22'b0000000000000001011101;//R
            7'h53: data = 22'b0000000000000000010101;//S
            7'h54: data = 22'b0000000000000000000111;//T
            7'h55: data = 22'b0000000000000001110101; //U
            7'h57: data = 22'b0000000000000111010101;//V
            7'h57: data = 22'b0000000000000111011101;//W
            7'h58: data = 22'b0000000000011101010111;//X
            7'h59: data = 22'b0000000001110111010111; //Y
            7'h5A: data = 22'b0000000000010101110111;//Z
            
            default: data = 22'b0;
        endcase
    end
endmodule

`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/06/2021 02:11:38 PM
// Design Name: 
// Module Name: Deco_4_16
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Deco_4_16(input [3:0] entrada, output reg [15:0] salida
    );
    
    always @(entrada)
        case (entrada)
            4'b0000 : salida <= 16'b0000000000000001;
            4'b0001 : salida <= 16'b0000000000000010;
            4'b0010 : salida <= 16'b0000000000000100;
            4'b0011 : salida <= 16'b0000000000001000;
            4'b0100 : salida <= 16'b0000000000010000;
            4'b0101 : salida <= 16'b0000000000100000;
            4'b0110 : salida <= 16'b0000000001000000;
            4'b0111 : salida <= 16'b0000000010000000;
            4'b1000 : salida <= 16'b0000000100000000;
            4'b1001 : salida <= 16'b0000001000000000;
            4'b1010 : salida <= 16'b0000010000000000;
            4'b1011 : salida <= 16'b0000100000000000;
            4'b1100 : salida <= 16'b0001000000000000;
            4'b1101 : salida <= 16'b0010000000000000;
            4'b1110 : salida <= 16'b0100000000000000;
            4'b1111 : salida <= 16'b1000000000000000;
            default : salida <= 16'b0000000000000000;
        endcase
        
endmodule
